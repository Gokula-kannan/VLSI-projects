module pearson(input [7:0] msg,output reg [7:0] hash);
 
reg [7:0] t [255:0];
reg [7:0] i;
reg go=0;
 
initial
begin
t[ 0 ] =  126 ;
t[ 1 ] =  44 ;
t[ 2 ] =  29 ;
t[ 3 ] =  8 ;
t[ 4 ] =  93 ;
t[ 5 ] =  66 ;
t[ 6 ] =  147 ;
t[ 7 ] =  74 ;
t[ 8 ] =  141 ;
t[ 9 ] =  52 ;
t[ 10 ] =  91 ;
t[ 11 ] =  201 ;
t[ 12 ] =  74 ;
t[ 13 ] =  119 ;
t[ 14 ] =  223 ;
t[ 15 ] =  174 ;
t[ 16 ] =  167 ;
t[ 17 ] =  231 ;
t[ 18 ] =  224 ;
t[ 19 ] =  109 ;
t[ 20 ] =  243 ;
t[ 21 ] =  49 ;
t[ 22 ] =  18 ;
t[ 23 ] =  54 ;
t[ 24 ] =  191 ;
t[ 25 ] =  225 ;
t[ 26 ] =  172 ;
t[ 27 ] =  99 ;
t[ 28 ] =  167 ;
t[ 29 ] =  2 ;
t[ 30 ] =  10 ;
t[ 31 ] =  245 ;
t[ 32 ] =  234 ;
t[ 33 ] =  243 ;
t[ 34 ] =  136 ;
t[ 35 ] =  84 ;
t[ 36 ] =  232 ;
t[ 37 ] =  40 ;
t[ 38 ] =  173 ;
t[ 39 ] =  234 ;
t[ 40 ] =  253 ;
t[ 41 ] =  76 ;
t[ 42 ] =  115 ;
t[ 43 ] =  134 ;
t[ 44 ] =  174 ;
t[ 45 ] =  160 ;
t[ 46 ] =  158 ;
t[ 47 ] =  152 ;
t[ 48 ] =  54 ;
t[ 49 ] =  4 ;
t[ 50 ] =  241 ;
t[ 51 ] =  193 ;
t[ 52 ] =  186 ;
t[ 53 ] =  67 ;
t[ 54 ] =  200 ;
t[ 55 ] =  216 ;
t[ 56 ] =  14 ;
t[ 57 ] =  247 ;
t[ 58 ] =  173 ;
t[ 59 ] =  203 ;
t[ 60 ] =  42 ;
t[ 61 ] =  52 ;
t[ 62 ] =  111 ;
t[ 63 ] =  74 ;
t[ 64 ] =  4 ;
t[ 65 ] =  50 ;
t[ 66 ] =  37 ;
t[ 67 ] =  68 ;
t[ 68 ] =  213 ;
t[ 69 ] =  188 ;
t[ 70 ] =  174 ;
t[ 71 ] =  134 ;
t[ 72 ] =  200 ;
t[ 73 ] =  28 ;
t[ 74 ] =  8 ;
t[ 75 ] =  11 ;
t[ 76 ] =  174 ;
t[ 77 ] =  182 ;
t[ 78 ] =  78 ;
t[ 79 ] =  33 ;
t[ 80 ] =  64 ;
t[ 81 ] =  138 ;
t[ 82 ] =  208 ;
t[ 83 ] =  208 ;
t[ 84 ] =  179 ;
t[ 85 ] =  31 ;
t[ 86 ] =  24 ;
t[ 87 ] =  232 ;
t[ 88 ] =  56 ;
t[ 89 ] =  14 ;
t[ 90 ] =  94 ;
t[ 91 ] =  186 ;
t[ 92 ] =  157 ;
t[ 93 ] =  54 ;
t[ 94 ] =  207 ;
t[ 95 ] =  224 ;
t[ 96 ] =  191 ;
t[ 97 ] =  28 ;
t[ 98 ] =  115 ;
t[ 99 ] =  253 ;
t[ 100 ] =  152 ;
t[ 101 ] =  130 ;
t[ 102 ] =  204 ;
t[ 103 ] =  15 ;
t[ 104 ] =  189 ;
t[ 105 ] =  155 ;
t[ 106 ] =  125 ;
t[ 107 ] =  238 ;
t[ 108 ] =  34 ;
t[ 109 ] =  251 ;
t[ 110 ] =  54 ;
t[ 111 ] =  241 ;
t[ 112 ] =  155 ;
t[ 113 ] =  96 ;
t[ 114 ] =  22 ;
t[ 115 ] =  177 ;
t[ 116 ] =  150 ;
t[ 117 ] =  14 ;
t[ 118 ] =  150 ;
t[ 119 ] =  62 ;
t[ 120 ] =  230 ;
t[ 121 ] =  91 ;
t[ 122 ] =  54 ;
t[ 123 ] =  46 ;
t[ 124 ] =  172 ;
t[ 125 ] =  212 ;
t[ 126 ] =  40 ;
t[ 127 ] =  191 ;
t[ 128 ] =  76 ;
t[ 129 ] =  111 ;
t[ 130 ] =  127 ;
t[ 131 ] =  217 ;
t[ 132 ] =  246 ;
t[ 133 ] =  145 ;
t[ 134 ] =  108 ;
t[ 135 ] =  157 ;
t[ 136 ] =  185 ;
t[ 137 ] =  205 ;
t[ 138 ] =  136 ;
t[ 139 ] =  228 ;
t[ 140 ] =  5 ;
t[ 141 ] =  159 ;
t[ 142 ] =  45 ;
t[ 143 ] =  47 ;
t[ 144 ] =  252 ;
t[ 145 ] =  174 ;
t[ 146 ] =  139 ;
t[ 147 ] =  237 ;
t[ 148 ] =  23 ;
t[ 149 ] =  89 ;
t[ 150 ] =  93 ;
t[ 151 ] =  91 ;
t[ 152 ] =  85 ;
t[ 153 ] =  142 ;
t[ 154 ] =  190 ;
t[ 155 ] =  88 ;
t[ 156 ] =  21 ;
t[ 157 ] =  223 ;
t[ 158 ] =  238 ;
t[ 159 ] =  165 ;
t[ 160 ] =  178 ;
t[ 161 ] =  199 ;
t[ 162 ] =  125 ;
t[ 163 ] =  117 ;
t[ 164 ] =  25 ;
t[ 165 ] =  136 ;
t[ 166 ] =  200 ;
t[ 167 ] =  62 ;
t[ 168 ] =  36 ;
t[ 169 ] =  144 ;
t[ 170 ] =  99 ;
t[ 171 ] =  251 ;
t[ 172 ] =  110 ;
t[ 173 ] =  40 ;
t[ 174 ] =  159 ;
t[ 175 ] =  184 ;
t[ 176 ] =  177 ;
t[ 177 ] =  167 ;
t[ 178 ] =  182 ;
t[ 179 ] =  231 ;
t[ 180 ] =  224 ;
t[ 181 ] =  116 ;
t[ 182 ] =  228 ;
t[ 183 ] =  81 ;
t[ 184 ] =  160 ;
t[ 185 ] =  240 ;
t[ 186 ] =  177 ;
t[ 187 ] =  24 ;
t[ 188 ] =  62 ;
t[ 189 ] =  22 ;
t[ 190 ] =  132 ;
t[ 191 ] =  157 ;
t[ 192 ] =  102 ;
t[ 193 ] =  55 ;
t[ 194 ] =  36 ;
t[ 195 ] =  16 ;
t[ 196 ] =  148 ;
t[ 197 ] =  16 ;
t[ 198 ] =  28 ;
t[ 199 ] =  1 ;
t[ 200 ] =  155 ;
t[ 201 ] =  184 ;
t[ 202 ] =  152 ;
t[ 203 ] =  22 ;
t[ 204 ] =  203 ;
t[ 205 ] =  40 ;
t[ 206 ] =  141 ;
t[ 207 ] =  213 ;
t[ 208 ] =  61 ;
t[ 209 ] =  43 ;
t[ 210 ] =  142 ;
t[ 211 ] =  125 ;
t[ 212 ] =  38 ;
t[ 213 ] =  50 ;
t[ 214 ] =  98 ;
t[ 215 ] =  248 ;
t[ 216 ] =  38 ;
t[ 217 ] =  153 ;
t[ 218 ] =  172 ;
t[ 219 ] =  20 ;
t[ 220 ] =  159 ;
t[ 221 ] =  10 ;
t[ 222 ] =  40 ;
t[ 223 ] =  189 ;
t[ 224 ] =  37 ;
t[ 225 ] =  37 ;
t[ 226 ] =  73 ;
t[ 227 ] =  91 ;
t[ 228 ] =  71 ;
t[ 229 ] =  194 ;
t[ 230 ] =  225 ;
t[ 231 ] =  8 ;
t[ 232 ] =  105 ;
t[ 233 ] =  7 ;
t[ 234 ] =  212 ;
t[ 235 ] =  225 ;
t[ 236 ] =  253 ;
t[ 237 ] =  32 ;
t[ 238 ] =  50 ;
t[ 239 ] =  84 ;
t[ 240 ] =  21 ;
t[ 241 ] =  40 ;
t[ 242 ] =  187 ;
t[ 243 ] =  239 ;
t[ 244 ] =  98 ;
t[ 245 ] =  103 ;
t[ 246 ] =  230 ;
t[ 247 ] =  97 ;
t[ 248 ] =  127 ;
t[ 249 ] =  4 ;
t[ 250 ] =  172 ;
t[ 251 ] =  150 ;
t[ 252 ] =  49 ;
t[ 253 ] =  231 ;
t[ 254 ] =  251 ;
t[ 255 ] =  120 ;
go = 1;
end
 
always@(go)
begin
    if(go)
     begin
    hash = 8'b00001000;
    for(i=0;i<8'b00001000;i=i+1)
    begin
      hash = t[hash ^ msg[i]];
    end
    end
end
 
 
 
endmodule
