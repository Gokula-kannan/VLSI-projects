
module xor_gate(input [7:0] in1,in2,output [7:0] out1);

assign out1 = in1 ^ in2;

endmodule
